library ieee;
use ieee.std_logic_1164.all;

-- This component will be used 16 times in total during the encryption and posterior decryption process.
-- It  includes expansion, sustitution and permutation processes of the Low and High part of the data input.
entity SBB is

	port (	R: in std_logic_vector(31 downto 0);	--low part of the input data
			L: in std_logic_vector(31 downto 0);	--high part of the input data
			key: in std_logic_vector(47 downto 0);	--encryption key, generated by the K_block
			R_1: out std_logic_vector(31 downto 0);	--low output part, wich is feed to a new SBB block, until the 16th iteration
			L_1: out std_logic_vector(31 downto 0));--high output part, wich is feed to a new SBB block, until the 16th iteration
end SBB;
				
	architecture beh of SBB is
	
		component EXOR is		--First process of the SBB. It includes an expansion from 32 to 48 bits and posterior XOR operation with encryption key
			
			port (key: in std_logic_vector(47 downto 0);	--encryption key, generated for the K_Block according to the number of iteration beeing exeuted
					R: in std_logic_vector(31 downto 0);	--this block only uses the low part of the data input
					ex_out: out std_logic_vector(47 downto 0));	--expanded output
		end component;			
	
		component S_Box is		--The sustitution box. It forms a 32 bit output from a 48 bit input, processing them onto 8 6 bits blocks, each of wich		
								--will feed a diferent S block that will replace them for 4 bits blocks.

			port (	data: in std_logic_vector(47 downto 0);
					s_data: out std_logic_vector(31 downto 0));
		end component;
		
		component P is			--The permutation box. This component accomodates the 32 input bits to form a diferent 32 bits output

			port (	px_in: in std_logic_vector(31 downto 0);
					px_out: out std_logic_vector(31 downto 0));
		end component;

		component OREX is		--This block produces the XOR operation between the 32 most significant bits of the input data and the output of the P block
			port ( 	X_in: in std_logic_vector (31 downto 0);
					L: in std_logic_vector (31 downto 0);
					X_out: out std_logic_vector (31 downto 0));
		end component;
		
		-- These signals are initianlized just for simulation purposes according to a combinational system. 
		signal ex_sb: std_logic_vector(47 downto 0):=(others=>'0');	-- employed to conect the expansion and sustitution blocks
		signal sb_pb: std_logic_vector(31 downto 0):=(others=>'0');	-- employed to conect the sustitution and permutation blocks
		signal s_px_out: std_logic_vector(31 downto 0):=(others=>'0');	--employed to conect the permutation and OREX blocks
		
		begin
			etable: EXOR port map (	R		=>	R,
											key	=>	key,
											ex_out=>	ex_sb);
			
			sbox: S_Box port map (	data	=>	ex_sb,
											s_data=>	sb_pb);
											
			pbox: P port map (	px_in		=>	sb_pb,
                               px_out	=>	s_px_out);
                        
			OR_Exclusive: OREX port map (X_in 	=> s_px_out,
												  L 		=> L,
												  X_out	=> R_1);
													  
									
	process (R)
			begin
				for i in R'range loop
					L_1(i)<= R(i);		-- This is done because the most significant output bits arte the less significant input bits without changes
				end loop;
		end process;
		end beh;
